




module byte_joining (
  input [7:0] Lane_0;
  input [7:0] Lane_1;
  input [7:0] Lane_2;
  input [7:0] Lane_3;
  input [1:0] ctr_3;
  output [7:0] out;

  );

endmodule //byte_joining
