module testbench ();

endmodule // testbench
