module wrr_cond();

endmodule