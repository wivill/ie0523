module qos_synth();

endmodule
